module motion_detect_top #(
    parameter DATA_WIDTH = 32,
    parameter FIFO_BUFFER_SIZE = 32
)
(
    input logic clock,
    input logic reset,
   
);

endmodule
